//-----------------------------------------------------------------------------
//
// Title       : Control Signal Translator Testbench
// Author      : vinod sake <vinosake@pdx.edu>
// Company     : Student
//
//-----------------------------------------------------------------------------
//
// File        : control_signal_translator_tb.sv
// Generated   : 27 Dec 2016
// Last Updated: 
//-----------------------------------------------------------------------------
//
// Description : Performing testing on signals generated by control signal 
//		 translator
//		 	
//-----------------------------------------------------------------------------
`include "constants.sv"

module control_signal_translator_tb();
	logic [4:0]state;	//state from control state machine module
	logic [15:0]opcode;	//16 bit opcode from Instruction register
	logic [2:0]alu_flags;	//ALU flags from ALU module
	
	logic gp_write;			//write value from register to databus
	logic gp_read;				//read value from databus into register	
	logic [2:0]gp_input_select;		//select register into which data is stored
	logic [2:0]gp_output_select;		//select register from which data is loaded into databus
	logic [2:0]gp_alu_output_select;	//select register from which data is loaded directly by ALU 

	logic [3:0]alu_operation;		//
	
	logic latch_alu;	//loads the ALU result into ALU Latch
	logic alu_store_high;	//write the high 8 bits of ALU into databus
	logic alu_store_low;	//write the low 8 bits of ALU into databus

	logic mar_load_high;	//Load high 8 bits of memory address into MAR
	logic mar_load_low; 	//Load low 8 bits of memory address into MAR
	
	logic ir_load_high;	//Load high 8 bits of instruction from databus 
	logic ir_load_low;	//Load low 8 bits of instruction from databus

	logic jr_load_high;	//Load high 8 bits of jump destination address from databus
	logic jr_load_low;	//Load low 8 bits of jump destination address from databus

	logic pc_increment;	//Increment the program counter
	logic pc_set;		//set the program counter from jump register

	logic mem_read;
	logic mem_write;

	logic t_gp_write;
	logic t_gp_read;
	logic t_gp_input_select;
	logic t_gp_output_select;
	logic t_gp_alu_output_select;
	logic t_alu_operation;
	logic t_latch_alu;
	logic t_alu_store_high;
	logic t_alu_store_low;
	logic t_mar_load_high;
	logic t_mar_load_low;
	logic t_ir_load_high;
	logic t_ir_load_low;
	logic t_jr_load_high;
	logic t_jr_load_low;
	logic t_pc_increment;
	logic t_pc_set ;
	logic t_mem_read;
	logic t_mem_write;

logic clock = 1'b0;
always #50 clock = ~clock;

control_signal_translator control_signal_translator_dut(
	.state(state),
	.opcode(opcode),
	.alu_flags(alu_flags),
	.gp_write(gp_write),
	.gp_read(gp_read),
	.gp_input_select(gp_input_select),
	.gp_output_select(gp_output_select),
	.gp_alu_output_select(gp_alu_output_select),
	.alu_operation(alu_operation),
	.latch_alu(latch_alu),
	.alu_store_high(alu_store_high),
	.alu_store_low(alu_store_low),
	.mar_load_high(mar_load_high),
	.mar_load_low(mar_load_low),
	.ir_load_high(ir_load_high),
	.ir_load_low(ir_load_low),
	.jr_load_high(jr_load_high),
	.jr_load_low(jr_load_low),
	.pc_increment(pc_increment),
	.pc_set(pc_set),
	.mem_read(mem_read),
	.mem_write(mem_write)
);

// Waveform log file and monitoring
initial begin
	$dumpfile("control_signal_translator.vcd");
	$dumpvars();
end

initial begin
	#200;
	//Reset
	state = `S_RESET;
	opcode = 16'h1234;
	zerosinals();
	checksignals(`__LINE__);
	#100;

	//Fetch 1
	state = `S_FETCH_1;
	opcode = 16'h08fe;
	zerosinals();
	t_ir_load_high = 1;
	t_pc_increment = 1;
	t_mem_read = 1;
	checksignals(`__LINE__);
	#100;

	//Fetch 2
	state = `S_FETCH_2;
	opcode = 16'h0000;
	zerosinals();
	t_ir_load_low = 1;
	t_pc_increment = 1;
	t_mem_read = 1;
	checksignals(`__LINE__);
	#100;

	//ALU operation with source register - first stage
	state = `S_ALU_OPERATION;
	opcode = 16'h08e4;
	zerosinals();
	t_gp_write = 1;
	t_latch_alu = 1;
	checksignals(`__LINE__);
	#100;

	//ALU operation with source register - second stage
	state = `S_STORE_RESULT_1;
	opcode = 16'h08e4;
	zerosinals();
	t_gp_read = 1;
	t_alu_store_low = 1;
	checksignals(`__LINE__);
	#100;

	//ALU operation with source register - third stage (only if operation is multiply)
	state = `S_STORE_RESULT_2;
	opcode = 16'h1ae4;
	zerosinals();
	t_gp_read = 1;
	t_alu_store_high = 1;
	checksignals(`__LINE__);
	#100;

	//ALU operation with source immediate & LOAD operation when opcode has source_immedite
	state = `S_FETCH_IMMEDIATE;
	opcode = 16'h24e4;
	zerosinals();
	t_gp_read = 1;
	t_pc_increment = 1;
	t_mem_read = 1;
	checksignals(`__LINE__);
	#100;

	//LOAD operation - first phase when opcode has source_register
	state = `S_COPY_REGISTER_1;
	opcode = 16'h81e0;
	zerosinals();
	t_gp_write = 1;
	checksignals(`__LINE__);
	#100;

	//LOAD operation - first phase when opcode has source_memory & STORE & MOVE operations
	state = `S_FETCH_ADDRESS_1;
	opcode = 16'h82e4;
	zerosinals();
	t_mar_load_high = 1;
	t_pc_increment = 1;
	t_mem_read = 1;
	checksignals(`__LINE__);
	#100;

	//LOAD operation - second phase when opcode has source_memory & STORE & MOVE operations
	state = `S_FETCH_ADDRESS_2;
	opcode = 16'h92e4;
	zerosinals();
	t_mar_load_low = 1;
	t_pc_increment = 1;
	t_mem_read = 1;
	checksignals(`__LINE__);
	#100;

	//LOAD operation - third phase when opcode has source_memory
	state = `S_FETCH_MEMORY;
	opcode = 16'h82e4;
	zerosinals();
	t_gp_read = 1;
	t_mem_read = 1;
	checksignals(`__LINE__);
	#100;

	//STORE operation - third phase
	state = `S_STORE_MEMORY;
	opcode = 16'h8ae4;
	zerosinals();
	t_gp_write = 1;
	t_mem_write = 1;
	checksignals(`__LINE__);
	#100;

	//MOVE operation - third phase
	state = `S_TEMP_FETCH;
	opcode = 16'h92e4;
	zerosinals();
	t_latch_alu = 1;
	t_mem_read = 1;
	checksignals(`__LINE__);
	#100;

	//MOVE operation - fourth phase
	state = `S_FETCH_ADDRESS_3;
	opcode = 16'h92e4;
	zerosinals();
	t_mar_load_high = 1;
	t_pc_increment = 1;
	t_mem_read = 1;
	checksignals(`__LINE__);
	#100;

	//MOVE operation - fifth phase
	state = `S_FETCH_ADDRESS_4;
	opcode = 16'h92e4;
	zerosinals();
	t_mar_load_low = 1;
	t_pc_increment = 1;
	t_mem_read = 1;
	checksignals(`__LINE__);
	#100;

	//MOVE operation - sixth phase
	state = `S_TEMP_STORE;
	opcode = 16'h92e4;
	zerosinals();
	t_alu_store_low = 1;
	t_mem_write = 1;
	checksignals(`__LINE__);
	#100;

	//Loading high Jump instruction
	state = `S_LOAD_JUMP_1;
	opcode = 16'h7800;
	zerosinals();
	t_jr_load_high = 1;
	t_pc_increment = 1;
	t_mem_read = 1;
	checksignals(`__LINE__);
	#100;

	//Loading low Jump instruction
	state = `S_LOAD_JUMP_2;
	opcode = 16'h7800;
	zerosinals();
	t_jr_load_low = 1;
	t_pc_increment = 1;
	t_mem_read = 1;
	checksignals(`__LINE__);
	#100;

	//Always Jump
	state = `S_EXECUTE_JUMP;
	opcode = 16'h7800;
	zerosinals();
	alu_flags = 3'b000;
	t_pc_set = 1;
	checksignals(`__LINE__);
	#100;

	//Jump if carry
	state = `S_EXECUTE_JUMP;
	opcode = 16'h7801;
	zerosinals();
	alu_flags = 3'b010;
	t_pc_set = 1;
	checksignals(`__LINE__);
	#100;

	//Jump if carry - Fails as carry flag is zero
	state = `S_EXECUTE_JUMP;
	opcode = 16'h7801;
	zerosinals();
	alu_flags = 3'b000;
	checksignals(`__LINE__);
	#100;

	//Jump if zero
	state = `S_EXECUTE_JUMP;
	opcode = 16'h7802;
	zerosinals();
	alu_flags = 3'b100;
	t_pc_set = 1;
	checksignals(`__LINE__);
	#100;

	//Jump if zero - Fails as zero flag is zero
	state = `S_EXECUTE_JUMP;
	opcode = 16'h7802;
	zerosinals();
	alu_flags = 3'b000;
	t_pc_set = 0;
	checksignals(`__LINE__);
	#100;

	//Jump if negitive
	state = `S_EXECUTE_JUMP;
	opcode = 16'h7803;
	zerosinals();
	alu_flags = 3'b001;
	t_pc_set = 1;
	checksignals(`__LINE__);
	#100;

	//Jump if negitive - Fails as neg flag is zero
	state = `S_EXECUTE_JUMP;
	opcode = 16'h7803;
	zerosinals();
	alu_flags = 3'b000;
	t_pc_set = 0;
	checksignals(`__LINE__);
	#100;

	//System Halt
	state = `S_HALT;
	opcode = 16'hf800;
	zerosinals();
	checksignals(`__LINE__);
	#100;

	//LOAD operation - second phase when opcode has source_register
	state = ` S_COPY_REGISTER_2;
	opcode = 16'h81e0;
	zerosinals();
	t_gp_read = 1;
	checksignals(`__LINE__);
end

task checksignals(input integer lineNum);
begin
	#50;
	if(gp_write === t_gp_write) begin
		$display("%3d - Test passed for gp_write", lineNum);
	end
	else begin
		$display("%3d - Test failed for gp_write, expected %h, got %h", lineNum, t_gp_write,gp_write);
	end
	if(gp_read === t_gp_read) begin
		$display("%3d - Test passed for gp_read", lineNum);
	end
	else begin
		$display("%3d - Test failed for gp_read, expected %h, got %h", lineNum, t_gp_read,gp_read);
	end
	if(latch_alu === t_latch_alu) begin
		$display("%3d - Test passed for latch_alu", lineNum);
	end
	else begin
		$display("%3d - Test failed for latch_alu, expected %h, got %h", lineNum, t_latch_alu,latch_alu);
	end
	if(alu_store_high === t_alu_store_high) begin
		$display("%3d - Test passed for alu_store_high", lineNum);
	end
	else begin
		$display("%3d - Test failed for alu_store_high, expected %h, got %h", lineNum, t_alu_store_high,alu_store_high);
	end
	if(alu_store_low === t_alu_store_low) begin
		$display("%3d - Test passed for alu_store_low", lineNum);
	end
	else begin
		$display("%3d - Test failed for alu_store_low, expected %h, got %h", lineNum, t_alu_store_low,alu_store_low);
	end
	if(mar_load_high === t_mar_load_high) begin
		$display("%3d - Test passed for mar_load_high", lineNum);
	end
	else begin
		$display("%3d - Test failed for mar_load_high, expected %h, got %h", lineNum, t_mar_load_high,mar_load_high);
	end
	if(mar_load_low === t_mar_load_low) begin
		$display("%3d - Test passed for mar_load_low", lineNum);
	end
	else begin
		$display("%3d - Test failed for mar_load_low, expected %h, got %h", lineNum, t_mar_load_low,mar_load_low);
	end
	if(ir_load_high === t_ir_load_high) begin
		$display("%3d - Test passed for ir_load_high", lineNum);
	end
	else begin
		$display("%3d - Test failed for ir_load_high, expected %h, got %h", lineNum, t_ir_load_high,ir_load_high);
	end
	if(ir_load_low === t_ir_load_low) begin
		$display("%3d - Test passed for ir_load_low", lineNum);
	end
	else begin
		$display("%3d - Test failed for ir_load_low, expected %h, got %h", lineNum, t_ir_load_low,ir_load_low);
	end
	if(jr_load_high === t_jr_load_high) begin
		$display("%3d - Test passed for jr_load_high", lineNum);
	end
	else begin
		$display("%3d - Test failed for jr_load_high, expected %h, got %h", lineNum, t_jr_load_high,jr_load_high);
	end
	if(jr_load_low === t_jr_load_low) begin
		$display("%3d - Test passed for jr_load_low", lineNum);
	end
	else begin
		$display("%3d - Test failed for jr_load_low, expected %h, got %h", lineNum, t_jr_load_low,jr_load_low);
	end
	if(pc_increment === t_pc_increment) begin
		$display("%3d - Test passed for pc_increment", lineNum);
	end
	else begin
		$display("%3d - Test failed for pc_increment, expected %h, got %h", lineNum, t_pc_increment,pc_increment);
	end
	if(pc_set === t_pc_set) begin
		$display("%3d - Test passed for pc_set", lineNum);
	end
	else begin
		$display("%3d - Test failed for pc_set, expected %h, got %h", lineNum, t_pc_set,pc_set);
	end
	if(mem_read === t_mem_read) begin
		$display("%3d - Test passed for mem_read", lineNum);
	end
	else begin
		$display("%3d - Test failed for mem_read, expected %h, got %h", lineNum, t_mem_read,mem_read);
	end
	if(mem_write === t_mem_write) begin
		$display("%3d - Test passed for mem_write", lineNum);
	end
	else begin
		$display("%3d - Test failed for mem_write, expected %h, got %h", lineNum, t_mem_write,mem_write);
	end
end
endtask

task zerosinals();
begin
	t_gp_write = 0;
	t_gp_read = 0;
	t_gp_input_select = 0;
	t_gp_output_select = 0;
	t_gp_alu_output_select = 0;
	t_alu_operation = 0;
	t_latch_alu = 0;
	t_alu_store_high = 0;
	t_alu_store_low = 0;
	t_mar_load_high = 0;
	t_mar_load_low = 0;
	t_ir_load_high = 0;
	t_ir_load_low = 0;
	t_jr_load_high = 0;
	t_jr_load_low = 0;
	t_pc_increment = 0;
	t_pc_set = 0;
	t_mem_read = 0;
	t_mem_write = 0;
end
endtask

endmodule 